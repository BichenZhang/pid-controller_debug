localparam NULL_SRC = -1;
localparam NULL_CHAN = -1;

localparam ADC_OS_INIT = 1;

localparam CHAN_SRC_SEL_INIT = NULL_SRC;

localparam OVR_OS_INIT = 0;

localparam PID_LOCK_EN_INIT = 0;
localparam PID_IGNORE_INIT = 0;
localparam PID_INV_ERROR_INIT = 0;
localparam PID_SETPOINT_INIT = 0;
localparam PID_P_COEF_INIT = 0;
localparam PID_I_COEF_INIT = 0;
localparam PID_D_COEF_INIT = 0;

localparam OPT_INIT_INIT = 0;
localparam OPT_MIN_INIT = 0;
localparam OPT_MAX_INIT = 0;
localparam OPT_MULT_INIT = 1;
localparam REP_RATE_MULT_INIT = 1;
localparam OPT_RS_INIT = 0;
localparam OPT_ADD_CHAN_INIT = NULL_CHAN;
//localparam REF_DDS_SEL_INIT = NULL_CHAN;
